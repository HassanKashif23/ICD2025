module test;
    bit clk,rst;


    axi4 stream
    (
        .
    )
endmodule





