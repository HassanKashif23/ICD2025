module parser(
    input logic clk,rst,

    packet.slave input_axi,
    packet.master output_axi
);

//Packet parser
    
endmodule