module parser #(
    parameter DATA_WIDTH = 128,
) (
    input logic clk,rst,
    input logic [DATA_WIDTH-1:0] data,
    output logic [DATA_WIDTH-1:0] parsed_data
);


    
endmodule